module lut_map_xor(
    input a, b,
    output y
);
    assign y = a ^ b;
endmodule