module lut_map_and(
    input a, b,
    output y
);
    assign y = a & b;
endmodule