module lut_map_not(
    input a,
    output y
);
    assign y = ~a;
endmodule